library verilog;
use verilog.vl_types.all;
entity tb_lru is
end tb_lru;
